module main

const(
	screen_size = 800
	cell_size = 20

	cell_amount = screen_size / cell_size

	// physics parameters
	influence_dist = 200
)