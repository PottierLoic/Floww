module main

import gx

const(
	screen_size = 800
	cell_size = 7
	background_color = gx.black

	cell_amount = screen_size / cell_size

	// physics parameters
	influence_dist = 200
)