module main

import gx

const (
	background_color = gx.black

	size = 800
	cell_size = 10
	cell_amount = size / cell_size

	iter = 10

)