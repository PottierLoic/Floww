module main

const (
	size = 256
)