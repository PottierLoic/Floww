module main

const (
	size = 256
	iter = 10
)